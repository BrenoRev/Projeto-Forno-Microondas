module t_input_control (
    
);